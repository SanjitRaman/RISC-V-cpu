module instr_mem #(
    parameter DATA_WIDTH = 32,
    parameter ADDRESS_WIDTH = 2
) (
   input logic clk,
   input logic [ADDRESS_WIDTH-1:0] a,
   output logic [DATA_WIDTH-1:0] rd
);
    
endmodule